module notgate(a, b);

 input a;
 output b;

 not(b,a);

endmodule